`default_nettype none

module Top(
  input logic clk100,
  input logic reset_n,

  
);

endmodule