// `default_nettype none

// module ProgramMemory(
//     output logic [3:0] out,
//     input logic [3:0] in,
//     input logic [7:0] addr,
//     input logic write
// );

//     logic [3:0] mem [0:255];

//     assign out = mem[addr];

//     always_ff @(posedge )

// endmodule

// module DataMemory(

// );

// endmodule